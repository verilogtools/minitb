// ----------------------------------------------------------------------------
// Environment package
// ----------------------------------------------------------------------------
package minitb_env;
  import uvm_pkg::*;
  `include "minitb_env_cfg.svh"
  `include "minitb_scoreboard.svh"
  `include "minitb_env.svh"
endpackage

