// ----------------------------------------------------------------------------
// Minitb types, parameters and helping functions package
// ----------------------------------------------------------------------------
package minitb;
 parameter int BusWidth = 32;
endpackage : minitb
