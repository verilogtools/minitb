// ----------------------------------------------------------------------------
// Data interface sequence library package
// ----------------------------------------------------------------------------
package data_seq_lib;
 import uvm_pkg::*;
 `include "data_sequence_item.svh"
 `include "data_workload_seq.svh"
endpackage
