// ----------------------------------------------------------------------------
// Minitb Virtual Sequencer lib package
// ----------------------------------------------------------------------------
package minitb_vseqr;
  import uvm_pkg::*;
  `include "minitb_vseqr.svh"
endpackage

