// ----------------------------------------------------------------------------
// Test library package
// ----------------------------------------------------------------------------
package minitb_test_lib;
  import uvm_pkg::*;
  `include "minitb_base_test.svh"
  `include "minitb_dummy_test.svh"
endpackage

