// ----------------------------------------------------------------------------
// Data agent package
// ----------------------------------------------------------------------------
package data_agent;
  import uvm_pkg::*;
  `include "data_agent_cfg.svh"
  `include "data_agent_monitor.svh"
  `include "data_agent_driver.svh"
  `include "data_agent.svh"
endpackage
