// ----------------------------------------------------------------------------
// Minitb sequence lib package
// ----------------------------------------------------------------------------
package minitb_seq_lib;
  import uvm_pkg::*;
  `include "minitb_vseqr.svh"
  `include "minitb_workload_vseq.svh"
endpackage

